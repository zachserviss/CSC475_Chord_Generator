BZh91AY&SYɿ �߀Px���g������P�rB�̀�	B�~���ꍵCF��4=Lj��A�101��&%2@�I�<��2   4�101��&$HML��OQ�e<�������I|Ї�I�J���$����$�F&� j}���bJѤ�b���aF�k��<ex����r�;h["Q#�)�|�bRzq1F6�H��O�b�k:uh�b�1&����xǠfD�����)^�3�@��HF�ǰ�W7���r� �z��Soh܃���'�
n^�ܗ����9ʺ�g ���Q������ Wf��]��#E��̤���J����o+9�+�%R0gL��QKS�&�W�6��toj��t��j�3u��.sbcx��l<��w�#�����լ�;ՉR�{��ĒI?*hӤRƘ�f��A�EƉ�y��11�Ȱ
�
�2����35OwH���S�6��Ea�Ɖ;Ǟ�߱΍e�d<X��|Q4`�����]�E�LZ����"nى�Ǆ�Y P�iI�����A���ɀj@lW�?r�!H+΢H�|��ٖ���Ѩ�NIzd9!�gDq�xf��ռy�	�7
��Z��/�r��*�)r�`��+Kе�!��� �����f�%VD�^�\��1�>����b5Ƀ�brȯY�ˊ���z�����Z���'���yKB�h	i
37#����x�"FC� V�#'�G9i�%5�3X�t��b�Ian\Kp	�X�Լ���l%�����҆�ZIj �z�F���n{�Q^vb���A����Գ��A��+�$�A'�3|�
B+���qÑb	db�jHܘ�5�Ӽs�/w�ah�l�eA;�P��ID3�@�'��fL�a�VMđy�!����}C�ZG��|=G�smWM �@8&4Ʒx#XH��Ȟ��{z.M�B��%V�H��ȼժ6+�ѳud*�k�0V)f,
��4 ���R��%���JU�E�m��XH(�:葆�6L\���i2v�b%�������m���_M�
?M�q� �`�/̊���H�
7�/�