BZh91AY&SY��H4 �߀Px���g������P�]��5��%?S���G�ɢ= �OPz���挘� ���F	� �� �M#���M@h3P ��� 挘� ���F	� �$ �S�F��yOҀ�A�jz����i'�B(�U� �~��%��16�HCP���M��sX4�L]�mI����2̔`\X�%o�u���ў�о��\���b�cY�F?�)�Ef��^u,TF����.~$��a(�ԯZY��H1�B0E\��z>gwu���0cy���-.�=�d�7����(�Q�;���
Xr�6��(�i��"�g��[�ٖ�LQA(ī��5*�kEYB3^E�&��8�7M���xx�����$�@��}�������tM��R;u��<5�R�{�?��t�C���ljbD��C)���Q\�1
;��BP	FHͽUz��ȭ�0����7�(��$�I�oU�>�?c��i8�.}��K��<(���!�b1�`�~4� J�JQ����b2tC�$�T����V#&#�P�z���,����$(G�J���1����^�HsD�����Z��I��ղ���8�Vqs#���-U�tdX�T�q0s�V����!�A�b��'h,
�*��r��VL3��^�dC��U��MZW�1^ d;�6���,TRJ����u�)b�D��	�Q�W%�j�L���aD��n;zT���a�7�^��d2B8�B�H���.������(�Ɓf"Υ�F/����9B2��t��ZQ��HXNjZ�c �2�+��a#��Q$�WF&�s���X�\F���&�A(&�uXw�2�q�X
��u`�ܑ�F|�9#"BV�6h��D���10�P3XŘ�5s��5��i��>�Ol�HbcLk�z3�$v~d�[Y��jh-�+�
�TJlI""�v�ުkY�}���*�3�/U)h*
)�v����jP���`5
L��^sP�|Z�����$J��H�y�&/S��L�H/�=
�d#n���|'�h�=�����8l�A���]����H�
���