BZh91AY&SY'� \߀Px���g������PXz6 �Ml$��i�e6���!��i��G�444d���`F�b0L�`�2jdM(�S���jyz���hѠѵ=OPѓ �`A��2`�I"{I�~$L�ڞSO"   =F(������$����(eX�H5<O��Id��0�#&k��㦁����%�#�r|�C9�s��V!�%�2|>&7���ی���У)���5&c+�nJ���<@���+Dx�}eW���R�0c�?uyy�̺��\붜I����;�O8)T�mf�0�2Ϫ�%�(jA���ɖS�_���si���kM��u61���m���=��.��N��9UE�Z̳窗6��W�j�����0�H1zC��X��X��������66�͑=�d}7˼�yld�>�g���+��?��Z�Clq��P9�i#k𺬃~Uz��2(&#�A��bٟ��`�br����w�		JQ���N`ͨ6�T("ۃ�2�d۵NbxKRs��~�<��b�@;����9C� ��`P�l��X��{�/���z��$�G#,���A׾�ms
Q��V޸���Ȏ�`�hRO 4�2�6dR'�������Zh-)2����3�1Q/	r�`�Ya�sV8�A<?�������4�d?P8 <5@؎��Ww���/ �[��}���T+J�-�5��lX�J�Q�(,&��{/��Q(��e�-52A�S�[�d\�F����U��5,�ʴ����ͱ�F��8`&z��D��H@���̄L
��bNI��E'm�cʬ���\D*�C���M�po�@G����5=�ˇ!Xq b���z#u�Ԗ��_�'rFA���u��)"Cu mL2a���&��}e�#ŅI�T`��"�A'���yY�.�E��gb�O�q�v,��d)�:ja�����B�- �h��4�X��xA'9��ff������H�%���EiY.2.�M�
�F㜍�
��׌6y�|�F5E��w$S�	�q9�