BZh91AY&SY�[Ԋ  _�Py���g߰����P�ck ��44kIP� ���aL���z���#��Q��Pz����2%j24�    �%4
b=@��MF ���a2dɑ��4�# C �DЀ4���zOTь�i��4�LEʤ7��@� `>� ������TD�H�{��_}�.$ \�w
6sk�$ۏ��>�W�<UեUUQUT�UUW�������|�r7�Gp?$%��=��BBRu��-�2;�� �5�r����VfE�1��$+�ډ5T�T�d�Ci{��e����1�p7UT��C�ݘ�i��2N ��������=@N�Wv�d��A�0�}��[krZ��A`������W@�$Lm0%�n"�X`x[c֜6!��[9&T�ǆ��͓�86��܊.A�K�]�M��E�1L(ĳ�ᢂ�/0�ide�##Zf'R�C�בO�S�IP���w˼�	�v5h1j&S�q�%z���81�5u
VZ����~X�u�q��m�A3�r�������Â(f�2�50���m�����@�� $6�"5�d�(�b�y^��\���G�ΊFaRD.��]#�@ @�% D(TNE�D��%�7�+�A�<�5�l�Q	d?>��D�@��=i5�4p�j�a(�?��ڸ��b�/���~����?8K&�\}%��ye�Z���TObI����s��<���&�=7���F �x��/��!̓�$��Q>A(�s)�r�jr�*4OO��t�ry�<K}�.Ie��e����!Qѳ��/���ێ��r�����Kmb+MJ����퇮��D����+w@
��!2�i|)ZW�ɬ��4'Ǵ�I��@�@�a��P���ѹ�%�M��"N|���3�s@��]��/�Wc@�%w�S����˕���0�@��]ċlG����,\�iP���� �S;�!:_nA=w����s�bh6��D�p|�D�:�c�tJ�2���F	��SaU��k7m��M�	����`T�i6�ڹ�؈� X�VmL��(��-,R�5�1��s R���]�Q�Nh��N<G�n��N��`��״�=����XD<ŌˁQ����@��(����k�s\�O�pB/��:DL����.�́��0E3u�F��F�G}c�`ag/��
���.jR�8IPtB�Q���5�B5⠂=��F �*29K|t�Hz%��K�*Z��}�p~�;�5+�v��^�[N[�0}
�r.Hy���ifР���L?�w$S�	�H�