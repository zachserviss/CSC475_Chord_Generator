BZh91AY&SYc�� �_�Px���g߰����`��>�  p0�F�T��$�y�L�Q�z�Bm4�j<������h6� �   4�ɓF�� �0F`j)��=6� �A��  2�12dф�14�&���
6"S�~�zOSA����E�J �\� �D�$�P��$߿���a"�.B
g�ɢ~2�$�d�G^���Q^��׋�������<�yT$���t�J�I)I(I$�$�$�J�d�I$�)$�X�JK32��h����Y�dir���TQ��ݝVxMLZ�Tgy�a.s*C�|��\�U��ig�3<d�ӳLS�[nE�Ld���߸�|>!���P� �e#,"�g�����%��ɑ!iNh$"��b}��_�6l�t$!0��xC�,�ހ)/[��]�6؂N� ;T�a����(i\y�#a�7�"q��q�E�w���o0�wR3��K7N�6�#��="�]p� E7M�09L"��1����Sϰ	h�H�`؇�,l���6�9��E[=a��źh�fM&��c&��lf&L�����a:̚��`!��v�*X@6�Qx���)L�f;��e0}]�\V�"�Iw+��n��T����Jt�k��bڎ�/fX��{!m�F��f=N����Z��;mr�3$n����D-S��pD �q���ww��c3oX!�Dv)�v`�X��c�K>m�̴;�=��Y�;2�K�5m���NA���ALTے"CL�}��F;�s����b�ט.Y�Z��l�v+�\��l�s�5�ie��О��g;T�o;K݂�W,����3��&�Yމ��*��BՈ�D9�)�e3�2�1��@�gW�Llǃ���A
+�UT��Q���*O���/2�M�b��Ķ�c�6*�R(��QΊ�/E�ґEQb��JQEX��,hj(��Qb�(�b�Tš��)EH�!Ȗq�����P����12Bf@!�R�N��������~�[��֚d��>^�ﶎR�yY�y����F�<�|u_�Q�N�i;��ĥ�����J��Y����� $/5oV����'�9@<��R��HB����Ykq\zE!~����Ҝy�5� ���K��rH�Qh�3!5���F2^�����G��'B;�[U�<�`��10���[�ѓ�tF�!��s��뀃n�Ү��Ş�.#��/��f5�`���� s�u�9�LĿ���@�n}A�%��b���]���<���ۣ�_�$H�͵,���)����ؤU�Whe��R�a�R�$�*�c5�?��ڧ[;:��C�ՈIu�!o���g�0=��#j��8t�F%Z	��S�ld�A��I	2'�3BDQX��P��6��mQo�h�J�7L"WÂ�f/�HP���=X�l6"t�-:In��RA���^Ґ�"Vh�Βh;\_0f�6���5����Ψ��HB��;���G4�-�'չ�W�,��$�ReU�	��Rs7988ԗ\�T��Ŗ�T����kf��R�R��ƩW�TC�31f2�B��ӕ���kJ��H�ϙ�,\�� 9x��*T�W(���#�j�v4�t�N�T����?��H�
b�w@