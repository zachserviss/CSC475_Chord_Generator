BZh91AY&SY#-�� �_�Py����߰����`�y�'Y� Z7��@P��M�z��h�M� 4S � 44=@��2�&���O(h0�  �0&&�	�&L�&	����JMDd      =@���S����=4 ��14�R	��!�驓Q�=ODh�������;
�rB(��+$��S��h��Vm>�U�����M�2I�u��S5�w�v��vvz�鉮��\{n��3df��7Y����nr6��>NNfff�\]�fF�ʹ��+}o�{�H(<���%*	~3�+3̕�s�����!�RS2)�ydJ�*�!Ed��z��[��T��yxP����.��z��"�]�n��0"���$�ؑ��m�d�LЩB���g�u�<�w$M�Z�0Y�%�	�p/e���{�K�MQ�,��`!�
A������"5���E5�hF�Tк�]�x�%
�L�v3��xf*f����ߔ�z�rv��e�H�S���b���:�x�f��,
�xR��I��h�P04�)�728S �͉�tN�%��4x�Q�n���&��u4�"�p@Fc�Sr<�gN&��"�B��d�bIۑ3Z�A�H�b�L夃=5����weO&��
�["�m�CpJ�!��y�T�4GZs��ˋ�t:s|��n���m��J:MJ1:;�;�Y�iA�V����M\�۵��0diq�[%��1��5m�"��v.�yr"[�utՇU������!r(�q+z�&cx��E;ks�zٚ=�c��:pR"������d�)Ngz����eP���Z�&��Ri�����,�fd�bfd�Rĥ�m��K2"�f	F*ŋ����mR�3%T
%�F�̸�����$6�H�^d4�	`ɫ;A���!�ȲasP�$3���^�窎,�E�bL�43uy���pi�,"w:���W��p����b�0�Gų$J�K�'��aE��@��FiKX���hޜ�Oy&�>
b;�g��h� �5hX��$� ~�lR�$Y AW� �=���9���"��K� !Y&)���I:Ҙza*$���a����޴��BID���;?N򅠯!�R� Hg�!R��<m�L�)��]q�p��1Q(�� E Ĵ9u-��|gx�B�/�/7�5'��qTҚ2I��K�y'bs���`k�@P����u���:����1<�A�j��Kn���azi$rЏf�b-Nh@�A	�q�,(r8v$v�J���6���M`gT�n*�O1&�?d�$<���&�l�C���IT*�,�i���JP�����%�')���XN���r�� ���&���I�"�񑨙�PǠ �1�Ê���u%Nk���"	p=�V���\s���[�A�D ��@�&��1��J� w��b���N�ҹ%���;���A.M �ǋFL.���@M��&�`|׆��/ɡ�Q¾ITL�a�H�}D�����>q�'d�5���< ��2���oĊ%t�0��w���H�
e�{�