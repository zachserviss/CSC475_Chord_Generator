BZh91AY&SY�i �߀Px����߰����P<����4dֺ4$��H��G�I�4z4h @�DP�O�I�dɁ d�F���  	L�&���h��@   "�jO54� �   D�j��i6��hFĀ�F� �]��ZF�P	@{��p\��P�V >Lr��@�d+������3�S9�0kj��Ϻ�ϡC*     I%�J��.���CI��[H"7�?(o-���T��	�q}��c�3#�,'�����9�Uk����$����s��m�]aT B^��m�\�������mQi�M�P�6�M��"Y��M����	<�)�CN��+8��(����13^TyUWfG�U�s��kdYh����`Q�wT���M�g9�B���&���&��h^�t��-N��,V^^��T[6h�˽J!�
=3R�2ۤ�w�.ln]�W3:nh��_W:�o)�]/�)7��IHIn��HDBb>��A�O	�bj��k2�JĩW�;��jytl�%��.&bbdp���J(�9������ꢺ0bw�#}	�	�{3DaH��W^������,�:�x��vu����	u��-����;��u��a�bd�&��d(�H��+d����0�3r\�����X�^�1W���� ��Z�%�D� Υ ��0��
	~���"�����$��W�:G4:"X�%��
�z5\���G��E
���4��}��WAK���[��V�D7�ebDr���L"��D��<�����;6��bg��i1��r�]�Rj�{�
����ǀ�M@*O��� �JY$�FgTT�2���EzD�Y�EC�R�Y���&�l|���n6��gq:���%M�3�kC�͜Ha��Б�Inܻ�4p����9B4�^���rȂ��B�sR��c x�A!��M�H)�	��q���s8���pmL�#|����;%@T�7\Z�L�J $�$7�趁ȴ�6���\s�����T�n4�>39���>�ɤj!��Y���J���a���ĘsR�������5���Y�
����$��׮6*5�5\�,-![1���UK�E>�j���䈈��
�P��
.{�`赜Z�
%Nj$_����"pZs��R�Ċ�ڮ �9��}�K�o��l�� �i�E���H�
��� 