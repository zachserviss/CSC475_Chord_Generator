BZh91AY&SY�<�� 4߀Px���g߰����P~we�pP:�Q?S���zS�Fj hh�� � �A��=$��A� h   4�5�h=@��@=@  i� s �	������`���`$HB2&S��4�A2 4�z��� ���@���b^ �k�𘕃H��sP���6�n!��P(O�����IP��!-��V\�/��椘�	B��V-�(Hy�	aj�q@D��D z{�c�ܵ��1闲����+~�Y���0�g�J. �YF��
�L(����*��h�K�8c���IC9N4�j��LZ�+!� ��Ӭ������S�D��$�oMAU;�%��u	+��3�ȓ��Lm��"�>�?z��\j�0fp{Yk\�C��=�8�!�La��J3���3S�v[��he�L[c�Llx Zt�*(����cLyO�fA���J�g}e��A_�"�R�K�f�.����qXM�ň�Vm�Qnz�n��gP'2)J�U��̧�;�2)�\��w�KX�jr�!�y`ƏR��K?�Lqq�P�9�+A���ay5B^~�|��Y�	\B�$����*ƒr(]j��S"_F�A�Х�r���^\��]ٕ���`��%�6��b�qr>Y5u#`ZVqb��-��O4�$�ba.�'P��0U�EL�\����PP�y�z.�9�L�0Ứ�;5���!q�A���й�gw!�[��h|i��lߤ.D��k�b�%]�F���I"�<.I��B�F�5eԛ����\�u^�E���@ՊU�65	���&�����dAn�G��ζ'�w�SI���7��F����"�(HKDQ 