BZh91AY&SY�fjL �_�Px����߰����Pgqiv.#F"R�II�zddL
i��L�@hh�C@�?@OJ�4      ="Ԛ��     �101��&"I4&�?)��zi�=4@0��5` ��P 7 L��'w��Y���dP����?�%��fEq�ݣg#aD��;qon'�sۡ��L�GO��I$�I$�$�$�I$�$�5�kR��.Ny򥬤�-�-�V��Y#$/ظ��f�9璹��q13�C�5�XAU3��R�b1��F#�J�b����1�ӟ�KRBL00����'Ө	ז�+A�� ���gg)��e9���fTÑMMK)te����0�
��D�.�-��e�@��Ć�Wot]��sIl(
6�k"�nj4�����xХ���d��'��G[�]5�Yͮ5��/��z�p�L���I����X��$QL��� ���5Pë�hi��و��).�3\Bū�
+V�,a�)���ͭ��cJM���P��!�0�����W�!\�
M��x�,�n��o=�}�ٴ/�4ۆ���UP��:��3d�WSh��̧���s���x�!!$�$�@�����=e/y�;"n��Tumi�w-I��b���i��.�T)i4�	p� �F���  �1   q��*�{��sK:^��}T@�.�p�� Ȥ�.uPv>�u4�%�7��~GӦ:&�~��Q��^���^��|��;�O�5ӂj�M��NY�FӰ��W�7yw<��m*Lq˨��^XD�K��� ���h�\Q{�B����=���p���4X������������}��!ټ�$�Q�	u��Nt��?�L����,��r��X�t����q0�?Kc��9�bQ��TTlW8#/���Z���������t�6����e�Kh����c�>g��8���FN��0�a�m�m���`ɵ�Ҭ�<k�7�3�dnk."[�L�I�+�4T��jX����!)��Z��$�A�N>x�ϙ�B�ݹs ȱ���[<�&��<�3a�Qx��ïn����&��E@��c��7̱D�!�|.$�Թ�r�d걓��fv��P�4��M�"-HK�9�@G�U���g����=�!�<����7����N���H�r?N��6��X��1���jqQw����a|���2��
��ve�h�zE��:�/yq�EJ�*)3�)��ѕӤ%D��U\5�!��6���ϳLs&y�+Kւ`�-v����ǎ+��l&�H�Ⱥ�׸0��dy�T11G��f6���502E8�G�]��BC���0