BZh91AY&SYE�F� [߀Px����߰����`�,�{�@ �n *��H$�F��E?!�54ɵ1=5= 4hz����	�R� 	�4    9�&& &#4���d�#���(�@ �4 �4 挘� ���F	� �"@��dS��i4���44�1z�΢O�!	!"�I$��?C���eX�H%I�a�{��_� .4��.��'���'e�՟&wh�~l5[
%)J2��&�m��m��m�M�-��m��6�|m��m��m����6ܶۖ���Ĳ�NC7���1���S��i�h�KJ84iL�$�L�ËOw�]�,TfҌ�ex2���yU�#g�-�c�!�0��f�N�'�����.�!&0c��<&� (1�涫��d�@��y;*�|�{Bw�wL�Sb�Z�教WW�bיUQs5C+�H��0��E��Q��h�;8(��Pe��z�����Ai�sU���$�jL'�Q�jQâ&��{`�6�hC��0�`Z�)IYRt�n��OMp�o���H*WYrg�9���:,�P8gA0�UT+%v2����ˡnc����:4G8�;���jD���'���������&!d�6,�Y+��tbq4A��O������z90���@���V����2+��9N���C�y���|r'W�5��*�� �b����^@p���,2A#"`At�T�5�R�A%$S*m�iKm"��B�ÞR��k�B�Fw�޼＝z�����z�VL��sY��u�6b7a���{������̠T"�
z�
Zy�Rť�#�y&��͋ Y�w̻Ԑʉ�ݨ��ǻ<P̎b�jD����$���,�{N��E+#7��|C�(��&11�D�k���X��x��^��;:��ok��� �m� 6�P�p�f�d]IP��.�A �Qĺ�@" @���`�"�bp��Sr��1�-ICZ����$6�Hmd��4�l�G��y{l��򳛉�4Ɏ�h?~'�}���g(���g�}��MX�M��h��Q1W����O1ZD�ǃ�s ��7�:�J��p���Yݮݡ���"�2� ;�F��f� _�D�	�'������Ȅ%]E�����61J�
����z��#�`��E�|V�_)wX��&����d�:1�Ď#70�H$u ��]"̉���xJ�������j5��hK"$rXqޚ�o9Ȼ���\��E�N�H�i�;T��I^�}5�\�Sƨ|C�x�̑[uU��ej��p�9CFGg1�p1��T�B��5\�c�N�~Kj�c8�[ �Kf��"��Zs�v{�\VK�5.�*�m$ZR�v��A$��� @�I���H�&V�8���\���C��aH;"Q�&
�e��Ad��*��E�0�&�Z,B��t߅DQ�L���w�p�^�V��a[���_x�c$e��5�Pm`͉�_j.B�;�-�ݞ)��;j��,ڪPt��GGDqUk�o9�tZ^E|�5���v
�c���B�D���P���r���{�"�$*�o�E
la��Ra��EAk���=���h�9�pe���l�IA���g���ܑN$h���