BZh91AY&SY�i� _�Px���g߰����P^u��[a	$E?E0��S�4�OS��z��`dz�s �	������`���`%4AS@�4��4���`&F F&&	�bi��! ��CI�&OMM2 M=M2]4=HJTH+AO��xHl	�-̆��p�H�i1t5
����5a��S��&@�T5��VI=���/���iX}iܙ"�g{��Z;���I�ӠW�!�G<�����K����&��Kf`'&Fg*ڱ�m���$
`t�Z��5�Iȅ%6
l�UXu�fAI���0��{��BUI$q̳�nWb��D�6����B�5(�����&!�1k$��k� !�5�{�ck�{�펻*�Y^[�����R�������;�<e�V�Eq��6��Yz�����yxl�N1���t��6�c�U�s�����ؠ6+��i�0�晴!�3i[�hB��G�������Z��=K��ql��E)]�p����r�@E;,��S�Q.4�J�������R����M*����`Ey��$���K��o���S���r�=Y��^�Ǚ�]$�>m�*K���2��U�X��Y�cX�𩆖H�C�Xt�5����;h{*%S�a�Y�Q�H�s�<���&&�Ā/$�M�*���h5�����_&�MU�h�N�$�ˀ�9�����>�Ś��:���H;y�J+&>4�DƵ��b�L�b�%]�F��Ã!4B��ooF�Fc�F
�
�4d���L��΍�iN��������)�yhM,��`��@^�����ND���Qy�z����9�����O~"�H�
M5� 