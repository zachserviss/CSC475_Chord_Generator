BZh91AY&SY�*� 
߀Py���g߰����`
���	��̑RV� �ZUR�Q)ꞌ��?<�eO�i���	�P�=(5=4JTi�i4ɂ0 !�@9�14L�2da0M4����%=$U       �A�ɓ&F�L�LDBh)��=Q��j<(�i �л01�YD**���@4*�}a+�L -4 R��0�$WLa��ta-
�k��^~}x����z��u��ܴXl����!�m�ke0�e��]]�M\����m7-��[-�w-��ܷm��c�h��{rݷ��oKE�/��;���d���(����5��r�B�B��JSJ�V��B��<��9q�j"��d�>T�i�Y���jS�c&U��0r.���ĕDP�l�f	�R��2�3Dݠ�вn��D�j���t�w���z��=1�P_���рf�T �'����	�Z�:��6��!J��o��9]����.�ˆ( a��#e8W(�cg~S:�ei\�ex��B������lË���G��8��	ʧe����9�v7��P!��ts���ǣ9�ș:0��Q�:9S�]��</KZ��ln+�+�Gka�0f-)@�R�MQ�8��!Uۡ��Pn�hkD�Jll�)��id3Pًق.������$WhPc�< ��c��C#g��o��>�Iv`��K�s�ܯP�%�$̺z d��qX:��/cvD��83��U�\�ʽ�9�aC�#,�#C,v�K�ep��CS[�3�wT��$G�M���� �^�EB���F�<�ֵ�#6փ�&��f*f̜̂q�5��gb�˺}�F
u9IH��ud1�\��prD�I�5g��$!c��q�J��ޜ�;,��M��NL�4(��b�����W�pNb�uޯ1:؋��B<��O��C�%@� P�$Q{�����ȡ J	���5q�͉���A�*���m��q!Q��fQ�/U�Sy�����î���<*�P��[٦�6c���e8�-
<?#Ǐ�q����;ToBk�k:*�A�:  ���u�
=�W8�,�&���g-�D0L�f�VZ����gqS��ٺ4V2�T��y��
��b�ZeQ�23��\� �&8�Y6\�Y�"���&b��̞���zwv{Yɘ�!"0`u8A�c0Md9�H�uAX��{"/, ͮߵ�c�����q�;��7�y� �OHZE|�UT���'�d<�8=��0�se���X�m��(��*�M"��ATU�@�(�*�H�Ѱ`���?�ى+(Њ"��#L�QDA	DE�JA�D�ADK��(����(��(�*b劢���*5�*���*�|Y'��HeX�aSE�����&0@�ѓY���tw�w�̺����a�Z����|vV�x:�(��<S�>����a���m�ͥ�K$�S�����̴y�}�.s��&�Z =�>�~��D�{�Cڅ�t �I	#�K\b�.�l�PI�ή,6?��� �װ��Fd����?>5����[ �I��}��Aq~�(Эk��~��b/,����/��F����HV��(�$44�Y��'��U�$~�ن�1��(6@$��A	��,���ڻ�mr�y� ��_+ں���U��oP@
NB�W!�w����T!<L��WT�����(��S+�=�!�}� ��s?(x�C�6���^�4f�
�@��z�/���FȤ�K^!���F�Pq5�P��A��Nm ���t7)B��rT'�!p�VB���!^�t�L���&Xb���
���E��� ���SIh�IΞ���\1�L�s�L�A��v�<C� _)�9ާN��fP���!��y�"�@�/S���W�2�7���P3�V
�$oede�FSȕ 15r\7YE���\��jz�ʨ V6��(��6��T^]�.-����X��wݎ�����w��й��)���>4ʹx�E\Ӗ8� �&%�j�?�w$S�	����