BZh91AY&SYҨT/ �_�Py���g߰����P��f��q��5�[��#Se�Tm)�"z�mG�I�@=M�=@�S
i<��h�=@     !"��$2h���  6�M0&&�	�&L�&	����=CI��F��=F���@���6�$�D@���`�@>~ce.�Q����j��n�f��0
�y\�{$A��]+؝�&\��Y"1���%�<w�0���c+geL�Z�k�l�4J׎�3s�rE77��T�̉�q��Ɂl$_w*�N(,YkL Y�^I$`�����9�qǎu�I�����4iJ�PW�ȯD!FA��,���b�%���f+C�#|���ph�]�-��q���1t��C�) њ$�V���,�ME�������Q�Qj�G��7�)k$�pAz���N4+��DaBMͫ&=:�_�������m��I������.�#��1WE��T�7T�x�*2=�*���� ����:�G�!le�w����-_<Dgk�[7Zc2�+�u�]>�v46Br��~f�h&��e?�
�xW.T���Z3ϥ[�;-XA��ż}dg��+�y��s�v��yAl{�X��D�@<��fk5���rp~�Y%����Z�B�� Ͱ"B�t�����̶�;���K1��sC�Pb�Q(_|���'�.`�pq��$��]%kl�6F��:M�R��s}�d��.̐�3m��+���N��fJ����,�Q��1��jt�bČbg�\��ʢ�e=�d��*����r\'�X��������o�h�ئ;��@��ߏ.Rƻ���g8�r��"�VҺ�r�HЮ�>������C��M�h�dė0��� h��9���r�^�B��23�i�K�U(��ld���%��P�	��$M2�c�F��-��L�dc�L��𪙓��f �@�g]��G3F�.��`��X��P����ң1�s��:�sZL�˔oP``Z�#ä�O2�	&Ґt�����%};~%F�fpi��@ӀU�D�nȒ  z�c����2�Vjt��HEpv�p�q�G^�Pj�&\�t�l����ԐQ(
w�
X��a��������9��c��.�#����e�ݍ�2�`�h֌�ܑN$4��