BZh91AY&SY 	�p  �_�Px����߰����Px�ӄ��6��I1�z�<�� bhA� �%*~I���(�    D���l�Oަ��@�i��ѓ �`A��2`�J!5�jF)�hz�	�@a_4�$�AD+@�����e l?]LP
Ƒ6�mC�U�MNDj��I��� �3����6D>�1���3h�d�2�mY�.'��� N���ak'��S�1�K��]{yr��K0���Cy[(���;@Őzo̺ot��W�ZB�%ã� ��{�!�\�kL���?��O/i*ʊg-)#},�����nRH;#���FS�����ء�}�5���UG�>�DҦ3I�}u�Y��b����3��=��g�0�_MOQ�YD�ۓ�e0<��S�;��w
G�p�p�,/\�j=���Y4��N9a�_�bHOZ{>��j;K�b�৕<�h|��"�����`P��tn� ����Usm���2�"A��O{��w�0�)�DkQQa[EY����3L�AZZĩeD��27aFP[U% ?�Cha��9V$O;dMJ1:>��Uȧ�x|��=���]U,����Y4f��
H�2q5q,Ƥ�C������4-ۖ����3��
\r��[QH�"8F����$Bd��C4���*�X2`9��%Y�șF����K��l���>⡀tG���b���x�!�.&����dV晷�"E�ӳ>(ӘX34�F�f�G'L�@��I���9e�����n�,��]p�d)��R�~p=��_��`��A�iA��q`�X.���b�@��׷]�W��fGɰ���~�a��!-�h/�E��w$S�	  �w 