BZh91AY&SY�,� �_�Py���g߰����`_-빺P �U�*�c���&&��CzS�SF�4��ڀ4hѦ�LJE  �    ���a2dɑ��4�# C ��2�P 4h�4�  h��T�@4��    	M	��%6������=&�&&� �h�� ?($�HL@����$���Ix2m&ЉI�a�~hp��#��d�H�,��[��s��$��v3��)�d�I �I$�I&	%�%��7�(�$�6������S,T��h���m,W#M7��2\�ao�U۴���
�,�����#�x�ۛ=EE)�eh�F;��gձ�*�f)�I"R,x�4`�}=�իi��5P$�d0ͽ�r��@�ɟM���s��	94Z���p�R����+���*E2R'SmB3�Ňf��p�(Z�&��[�t5�k��IJ+�Ό��d
U�Y�t�3R�k�\�j�Jz�
��F�q&q�&�!D�t�^�\l�qpÌN�&Ia5i����kv��5wP/' ]�-0�`��F:��UC��3���Ef�%�x�\$l�2�*YB3�pȴ�7U<��Z�0�N���%��##�C��L��������i�P�L�D�� �\�଩Q-wI)���ڷ2��X�"���[��^�I|ksh���-�O?�8��Ey��������?�x"�*�h�{�'z�M8�
��aE���d�uTUTjbEUEQEdeEUURFUUEY�E)L�$GW�֣[��/�`�C,w#�� ��Ս[t����t��}��ڸ��q���|�;tL�
uu��y���E�)�?ؿ/�T���I�n;��Y�	�]O*�q-+T��P��9��z���*��� 8��\k �*��9üc�Z�����IG�\<-�4�X/��IxR�`I6I�4�G-~����:�L�t#v9���ZmV��=�k��^�j�$o�AM1h	ԁ�NwE,�D�v�R#�aM��ѭLELD64�lr�U��j���ẽ0=6h�*�����{7��y�BJZ\�F�Q�=!��@�z�Q$8Yo�+[ժ�eƥB�T,+ļ6���*�N���zȵ0�b�1�I*fq�{pLV�0H4�Kf+�E����[=��R�+RD���x��TX��A�*����	w�$P�:��H̉��7��	�bMЕLpb*�.N  ���2;CɒD�@;e2�j�uM�a<\V.r��2���H�W��L�����^�	��5���eaBORX1������6:wa=�+8LrA�6L.���������v�V��ʲ��F�E�
��I�iH$��-�N�����Rf$Ã=�֌���tb< ��U��fax�b<qZK~#�,�L#�4�wQkh�4)��������0`�����"�(H~��h�