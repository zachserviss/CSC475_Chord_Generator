BZh91AY&SY��� �_�Py���g߰����`�," �jdѡ�$�2��'�Sd�M�h� =@4d�������@  ���&L�20�&�db``�����d a@ ���&L�20�&�db``(�)�jFJ~��� ��p
C��� ��?��@�/����B�a*��)���E�� 8�&3P��&	��b,�u�n��&�i���RI,E$�J�d�IRI�I)I(I%	$�$�)M�	V����Q���C�~��Op�8��<�,)��&b!��������jdSә$���'�'��߿����3?V]%"#�1C�7���x���ĕ���j���@�%=�$�hG7'Ӹ�R_�s�ҪH�!�n����*��,��+�7C�q�D��7���SҖ���-˫,KWf}�Wr�2����S4�V >�'��s�,>�X_��g02l�fr%7J����,m8]�;L���g �4Ȁ���T���e�1���0ڗ��S�Z� a%�6�sZ�͐�m��Y�8Z��鱫]	��|z��#��c4`���'1��h&[��h7W@�ú���Uw-�ȗ��^E�(�=8�gDLr�K�
��C���4��f�D[H�꺭�V-��w��M՜�Ɓ�Ox�ț�aGNEL�rr����/�,�e���3����ˁ�9�rY��〉��C�rXr����Yˇ�����	Af��^��%��!:��AÜ&v#��j����)�QWmQTD�!�pv^����l�;-j�x��T�a�i"����Lmt��ZUUUTd��*���*����"و�**"�b�����`�**����JeЪ�O����;涯�Q2k�l<-B��mk�K�Ϧy]\�妯'�V���$�u�tG��ۯU_�Ϗ���>s�I�OX7Q�o)N�f���ܔ���6�N�T�O��g4��������;���6E���p�U��_x�8��'F���~��1v(��r�}�%�,�4�l�~�8�*5�x��e)��b�⏀��s8j5��h��h�?�}�s���䒊�B��P�A��&������V���l�C`�C��T`�E ++�ß��%��.��"Nl�a�3�s@��]��۶�K@��^"�b��Jk��>�r7"q{r݁3U��Pd2��;u�Ij��PJ�ܡ	�}y��+}��s����A6�_5Mg)�9�h�Y��	�f-�Uz8mf�RB)��8J�D������-T]I~(؃"��[��*�BVC�v�ְ�by��n��أ5�8�v��}]L��Zw__i�7��ΟEr
��ʔ��W��O�8�;�'��z��$ء����;�	�T��.�́���L��`���e�gq88���,�&��VN�f���%�
�����EP��дd�^D6�Y)��9��)���Ve�X]�����r�Rb��f�\2��dv�(�b}Zݘ��#\~��.�p�!!S