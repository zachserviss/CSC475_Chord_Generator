BZh91AY&SYu� _�Py���g߰����`_,l� ^.%

D�$5=S�O�Jy=(=G���@4��4�T�D�%B�OPh    `LM&L�LM2100�U?T�i�@ L�@ �A�ɓ&F�L�LD����@��2`I��l��A�'��h@>@BI����1 $�q�}Y6�hG� 5=?����I� �aoi�A�'`�-���sj��\6S�[*�R��)]������www���������www��t'(2_��G��Y"���R�	�l��H(MivE�DTE0㝯t
r���������=/��©��d���3x�YB�g�ޖE[��@(�S `Zi�/�j�p�� 0�a��c>��}�l�јE�xA��7�R��,u�9�
�VF��TI��z�g)�u�D�B���`����ͩ�>��!�IRy�E��jV �G\�A��D�G4)���\",S|�!����&A6���]:�Q�����j�n\���֛�l�n �˷3X�X�oa�1)Cc1�B@����dkV٨���森�T�* M�w���QK�U��1��OLF�d�[Bҽ(���m	�_'WS\�U2&HoL_6�:�S��qtƙ՜���ky�#����7��������lA!D�o���`����sU|�S���kcf����?���-�V\�r�e=�Rd\�rIUU'"��Bp&2��Ñ@���"+ �8B
�L�"6H�e�W�0j�B!��j�Y���̪e��,�_��5H�][��_j�@ˮ�>4�9���OM���@��C���ν�|J��Օ9K���v� �j���p[��T{�V\��Bo�Y�W�;>�@xbF���^h�g�8$(G�ω}e�ܐ=R�}w�4:	�fT��rT�!޺!����c�$���m�Y��h�ی�r�)#��{���8bFMr&�
�0i��"Q-�2U���+��`5���X�C@�ږJ��V��5���{/�n,SP�I�]��>]U�j�\��
�k��K�)���	ŒpW6�o"X��
K�fm댷9� J���W�@�*J�>�l�&��6 OJ�@ѓ�l:��Ί��ň���5��ޥ�d�@��I ��H��2$�4�ZH���n*��T���b��� �u*bM�� T�.���Ѡ v���͉z3������`�9���=�q��˗�}A��u�����1ڮ&��@tZ�?��  �:���XZ]h4�L�AV�92!;��E����ad�e�)���5.��� WY���9����Rfe�-U���� ��S�'V�^aw'���d�V2)+���{���m&��������6�+�y��H�
��  