BZh91AY&SYO� ߀Px���g߰����PL�����	$�S�4&hO�1��P�i120	����L&i��S$&�����di���j s �	������`���`$�Dbd	�OI�6��   z�eCaBNI= �	6�����%��2�vQ0�A��"94�`�w�����8)(���<�%�K��O����g�V5(X��8@�j�\Y�H�n"����H�&t��<�i(:i���L4d�~: �XE·(���薒었`90�h�7|Õ�\��Aб��Ɗ3sxq��S$�$$��H�v׊9�RhR6V�+���V-d����.��p��TуQUF桉Fu�������s�_Nn>�t�O'W�D��C��8���.�v��l�\ř�pi�E�ѹ!9��B��:�R����ȇ}�f��Y/5D�@���i<V���*����#B#m∄>���M�p�Tk|m�x��<[�Z:�p��j�d��(fi���R?[ITXP��0B�:�AX�{��Ȩ���#��j�3�Aojۮ^5~#��0T�/n�R\�s�1^� ���=�2�ʲ�R{UJ8iC&��aj1��]��T��!AL+�E����m{�`~���!Y���Dh�dly,ڋ�a�/.�����7���`�Ǚ8t��6'g(�t�.dy��4�"7bF��-|�\�&��)�������=��
Re�T���kS@&���W0��E1��hk+
� ������-c["(`��PU~D7��Z6�T��`�p���e�^O�s,l�kp�rE8P�O�