BZh91AY&SY�k�� _�Px���g߰����PVy����n���MS�<�ڧ��Q�zi���dѡ�D����M����  �  @	M��)����G�@0M1�s �	������`���`$PSh#&E<� ���� �U!�BP��A4$�;H>�1,���R�=%������&tSYg�l�ɲ�vi�T5��M�n���c_P�k��k�$�I{�r���`H���vR)��R���̪�.5��Q�Oo@�#G�'��^dO��QJ�o��E3�'�e�D�<j���a0�B�I�޹Nv^2BVI$q�:gmƝ#Љ%�ґ�B*����^S jD2gW�Q��U6��BM�z;�_�w�xK^ǃF�lM�)�f؊#R<��;֐Z��>�5�v#���2�*r�!&RӸ$���!]x�a��Ў�=�cȬ4�f
!VJD�'���3R?�>y�¤3-����LL"�k\��#��'Q��[��m;_��W��{&�j�0��dɜ�d.���N����֦K��+�� � �$Pp�V!���E6qS Ԫ�nʏ�h�#Ƞ������"w[�3S�f�F���^�
���؆��X�{�1m2��b��U���"lW�E����;㜈&&���L��Uu�ycll�F��U�5N��!v���)���*��V�N�0���3#D��(%2r���o9�lT��7�5����4��L[��|$�4A�ay�t-�.Rf۰*�+�u��1��ҹN��=6��� ��uƠ���$0�l�Y�t?A��GZ����z]���Z�?�-6,����)�s^�