BZh91AY&SY8�6 ._�Px���g߰����P^r�p�B�0�)4i�g���4�!�50�4!@z� h    4����2Pd@4  i�)G�A�C ���  	L�L��I�2i�d  �Mh��{D�(	}��ؗp��k����v�Z4��t5
�k���\�    !8{H�<�Ư��ꇂ�B���F��eD�n�m}��Qe��^�	�%�8��.0`a�C�W���$ S��! �Lqz�3^xa+�E�����Ä!�%�T@Li�z^�pp�qj4�@`�6��P��cIL�B�L�-n�B`���w�U�ͪR��C�1*3)+��"�
S8FF�şB0��	DQT�DLAVRP�a�T��
H�;<�	��ⲋUl�U���G�Pq�1;���数������()e�0��NjKTx� � "!CMd��p�,I�)�UiI�~�I�i���%���SX�I�hM��� B��S34�4�#z�`�	�Xm��7�{撮RJ�e��s�n�`գ^ʄ�n��<��/=6���7����adc��*cr�9;
L�)^r�BB֨���ks{�D|l!|��'JRz��'��	.����p�}]B�!oES\	�f�*�1�Q����G��	̊R˪͇*\���N�e��ƃh�7J	o���E��E���+y����	�$��b�>c�XݳPci�M@P�?J>��*�Rȅ�D��~<��UL�A慲R҉d"(��V��L��ɱ�^�U����C�m5�\|�0����_�ʊ�0,3(ő$a9��2XB&�Ȁ$�H)!��~�����q��Eb��(	B�o�oy�j�I
�ðc�V�W,'�-��Zdh�f3��T�"�PQ���� �!�!P/�n�l�mĒ!@�/3�6*�3^{4� ,�ٍ0�*�[t�*Zo(7o/�B5�Y`S�xК[�45iC� �f+�k��3/�umU�T��A/���H�
Ն�