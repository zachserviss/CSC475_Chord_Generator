BZh91AY&SY��JH �_�Px���g߰����Py��s�c�h
�0�������jzi2=yG��L�D4hd4��% 2i�� 2@ $$�&D�4�@  �@9�&L�0�&&��!�0# ��I�d���)�d�T FM,�|@!%�	`I$�?�K�̘�P a�9,�,ƒ���A���O曺��ow�O�6w1wwuwf�����ɛ3�1��2��tg��vSUj��[P�6�˙t���I������u'kt~uځ����/�+y:�5����,�e  -����'DY^mh��<nL@��@�Z������5⃫�l�p�I�5RY�<&���XGm�e��l�Rj�v��0�ͱj�،�L�WS��i/UR�x�WŜ45�|ʈ�[)gD7���A%'j��>Lɽ	�P����GK�y�����2аaʠ\!�",�%�B����aȤ����ͻI��2�(q�u,M*�p����dպ�Kd���Ku��05�Ê�eXbf�m��![���7�A����`Ђ?�y/Q	|���M��JU?J��ꩍ��;:�mS#ln��cc�����jI$�J16�s2�])i�ի�3k���6��I��5��O�y�x؟[f~�T(�5E�m�p����E�z:�%�tT��]��B%���a��I�Z&U� /�h*�it�J_Ab\Ɇ�����805����@tX�=�v�HW�D��Q�'��w%�f\ >�AO�_�c�F��A��e�k�j��F2^�*��n#�ށ'a��ݩW#�2��u**G&X�M��$�1SH:-%Ev ��Lb�D�M��%B�|=n10��iU�Ms�U�9h��������:�n����ZY�����ڠN�BC>h�E����3��J��4~{�.4ܬX�Fc�u�`�nȡ� ����|��0~�I���p�C�&M [�>k���iq����gEy�ʣQF�i ce�v��A$$�� �Q���"��/��9��������a�.S,��5T�>��S̄@�M$`�F1a�]yH�8�CfJ�@��!b�xy-
�.)�Zu�x�,`�9�x�1s�@�4I��=�8�q��zh/*,u���J��D��TkM�x,+"�����U9�5_����ʈw``,B�m(���_-���P�FF�r��Q�I�^��pZ�����uo��)F��4T�3��F�Ԉ8X4�����"�(HGR�$ 