BZh91AY&SYw��x �߀Px����߰����`{pl��{��iEQJI�z��ZjHH�e<�OL��hP�i�M�44hz����茟�R�@d �i�  j��#U@b�22i�@��I��	Q��� 44  4m@hɉ�	���0 �`�0�I���23M4CL�  ѣNj���"
Z���
ʯ��;�i��@�����y0�?�I	��k1aF��\/|y�2�徧*ֵ�j    8       @        �4       �    �    @    a '��(���TF/Q~Z������XHN����
�B�i$�g\"E�*�Q�9JT�54�l�σ�CҼ�&Hf�����9�6W�	��r���@�]i��&g�p1>�3j9����E���>:O��K��oL4��ֵ�kZ֕���ƭ\�-����
@��Q� �2g�%	"F��ID�q�I�C�I�F��
�]1�Qȁ&(�N!*4�I��3�"g�X�4Z�b���6�� �b&B�y4f�w�tx�W#�[� ��?�g�c��Uф���D�^��Nt.��������(�U�7{��s�i=>1���8�Β,窝URtɲ櫤����VZo�;q��`���Nw�T��붮u�[�SN��8�wwV[���8k�[)�0��i�p���T�Oma���e8�V�]L.���P�m#9��ٶ�l��G^��m��O��L�&�h��E(o�]r��֡Օ��oUhe���}^.���dQ���"9��έ��tK!���N�:s/��<�ZGL�l���wn54�c���m��{�f�� �\�-ekP�bs�3��|\Z��l�w��u"���@<�ىԥW���o5a[y��en�Wɺ�[��,����m��tG���Q6�&Ei�Pə�|�|$Q�pPԎ�A�S=�k�G�w����6���.*�fw{�'8�N+v�ţD�&��`6�m��Z�r�
w
%=]iS��p�mK6����u��%\�l|�V�5:B�fcZ���M2�*�w�����Վ���%��@�HH�ҪORu��%�x�������ޕ�X�T�
���!��y�Y]9��0���W[�����ü�1�۰ zn����R�:|������q
��m�(�$�&RzI�93k��s�����9�Qj6D�1���(7����� ݯ`M����B^�$r	h�z�~��{��'T��y��:}�J�Z�"�)��ޥd�K[�����R��1aX��u�oI��|�  �D����37e>��(W/9\����/&��Zw]\\a>�cl��`�{�o^����/x���;�������UA!	(��ϳ<EI��?��������f[n΅QEEQE��TUTv�U5H,��R,H��Jan*��,�%�P
EUb��J�,QAb�X��e1bŊ,Qb�cB�,Qb��,X�b�#X�b�"*��QTQQEQV.�����s]3<PP����dĐ�$�ڵ�B���{)?��[���g��Ni�u�O��"���ߤ�[���q?:�'����������[3b���5fH�����/"Xs��v�30*g�~����������ޚ�_�(Hx+L_��8�����F���Ǌ��۠�k��DH�"�&x�/m̗�R4n��m����ŋ	�-���ۆ�-���I��O�;}���p�S	;�'�Ba!$(�T!��6�4�ur��K���/��bC�
���"�M\2L�>���������#�g%42"-5(xӊ^�G�y]4������V/�A��7Á[օr�$o@��>�s�Q�T��G{8oC������]�4`��o�����M�y�zIXCAA��h��	'=;�I(�Y��w�!�����>�����a�oh�d�lD�se�_��"�Pېᩯ 1�Қ�E�Zr�ѯp�k1��������������A�k0������OV��g�rX",l �md��ԛ�"�H����;u���
��%u�6�%�Q ��3���L��_H��%+��v	V�M��&fu`��
�9m�.�9I�ҁU��T��1��g��& �t�0r�қ�������Cr��S�:ᬊ�"툧�.�p� �n�