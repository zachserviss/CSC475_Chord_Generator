BZh91AY&SY���+ �_�Px���g߰����P�g��Hӭ	BJy����2�d��COQ�@d ��)�AA�     $%4�jG���L��� ��Ph9�&L�0�&&��!�0# �A	��$���I螦�M4  3� ��`�DI=�m/�,�؂�5}�����!d4�,^6�Ń�2�Jm�ŏ%U��Zՠ�c��oepH��dDn����FfW�b�Ya>؏�EEǠ|�q$DR���U��[��\\��Ͷ�-L
J "Q�-T"�Eg����L`��V����EkA�L<����֗��4��W�rcr���2��n�����9W��$�{R�ȩ�V�D�����eAǌ*19�%ģE�zV+�T��9�ib�/ѬƘȤ�V�����}����-���~-ʹ��5�U���)�ZFsI��K���`�0;:tFI���͖3����V�hk��f�UR
�����Z�Ǡ|�C����NtX�Mb>�?_�@��XR+�}�D��ZQwt�n���ă�G�n��88�~�62���K�(&ğMTg����Y#��آ�f���Z�A}�)�t�_��j �>��:q����
/�̝S�ߺ�r�=r	<	�c�Z�N-FN�K�QR:~���f��8������� 0i��T�F$__?"����wK��x7\$�B�X�XU�^� ��g,�jJ����sK�7�B�$dCTm�Z͝Dy�� *M#3���K���e؇%вՠ�	��C1�^���#T��Ɔ��B�v��Fg��xާ#	�C)Z2h/"+�%ƙ	����̀��Q��;�2�Q �x�XD�,�W�8�%/�S2yb�QX7l���O�b~�B;��P1������XW�ӣ�7�ٖ��b|���f���I,H'�ȘŻ���DI��z�Xp�h(歸*l�P<Y���Ӧ����k�]dEe�H�ԒB �)\ȂJ�eelv���S	ٖ�X���UQ�P	�E5�qb�P�"@�	)�Y�R�B��0S�T>K�"��C*�Y�60iʊ���H�
��`