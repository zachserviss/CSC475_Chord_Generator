BZh91AY&SY�!9 D_�Px���g߰����P�d.��(�'�����h���dɓ@���Q���� 2i�     ��&��h d�  �L9�&L�0�&&��!�0# �44�M5CBjz���d��Q�&Lh�'�I$�
������9_FU���&�����J�b�bvRUd�����~�暑W-k�    T 
R��  � ��UO�ЖS,SD��q�1��E������D���-��i��c���Fqe#��c�f��(��j�K%��� E�5JB2EK���jdww^��1����8�3ѧJ�nWAglڑ$MFLN"o9��V򛪚
v�k�a�[k�
Q�{��[^پ[��+#�(%�"{�zF�4��f5[�U��\�oj�BLL��1<B��*�T*�j�-+�kZ��X�m����9�'eN���Ģ��)4�*j1���f�g+9�\�j0�u`�8��b�}�
F�n�E��s��oW����ڧ֎:�^
8���	[��;�S����]���w�P�� D$����u������n&�Eµ�guT�v��g�� �54ڔKL�@ �p� &��!�&(i��b4بH�eO,ecXɫ����v�f��l mAE��eO�z&q�'�F�g�eEH�36������!����*������0�R*:��n�F���F�[�0��J@`����xf���Ay OT�^*��X�����p`�B����,�����B<��]��|�k���*�R���kP�Db*(_;+�#%��e��q�	:����V�:5�����~�x����tdBA���hD���tẺ���h(X2GϤ��I�k���Y��Ɓ9Ķ&��0-�j^�,��ŁeE�\S��U:�R�h9�$5����6т�1�� �B*梑娣S�iP�jB��~Ki~��)15��r�k︛�w3��28�I-���G�m:�0�uX���Yh5�QN���#�A�'	(	?<�D��eo�3�]DF ^�Z�t�D�S,��z�*��;/�5�0ٌh��4
X�ߓ&r�y�B�������W��=���G��|:�i�ΰ�> i�\<� Z�'��S�&	��;*��6U(9�� �X�T���C�v��3�#앹�$��F?� Wa$DFyC!K8ʇ6�n�-g�"�
�]�H��i͋�A�P�At�����G&�Zd�<͊�e���l�A��H�J-���)�	Ș