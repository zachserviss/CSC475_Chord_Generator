BZh91AY&SY��$ ߀Px���g߰����P^t��Um�J"j�H�<�?Jz�D�#��L@4h� 9�L�����a0CLM0��h�z��@ ���  �0# #	��14�H��Oi�x���a   ����BP��Aj}?�lK���Y����EF�c��`X�_a���Ɏ7�sMz9W�N�q
m�Y�Ϭ��L��k� �w��f����K$��G�?���Ӌc�/e7��Th�B���TD��fZ5�¤� 5YT�,qˁ�V���kz8k�761��km�dt�¹!�42rۈw\P:uC*�S5\�B��eD&���Hj�xL4�6�}Q?��=����/�m���p�>�b!}�.�Rʧ�u�j���u����CR�0yM��ǀI)I�)ÆԷ9��HG�}�+*����<�0��D#��}����|�-	���+��TؘF9ؽ��^`NdR��f㎅>�C "��˱�崁��4�ʌ�����u�J^bU���26*�qb]�CD�ȑ��eC�,M�
��&1�Ux]�@��KH&�7��Qy�Is6�ǶW�Y�fuɱ�ZfItTT���
	yQ0V���;������1dI�y'�X���]��&�di��J����W
3)P�D�S
ܴ�,'~1�_�%��vr0�I�F��+��C�M=�Ns���)�p�ג$Y3t�	+jl�lĒ!@�3�5*3F�X+ ,�Ս0��d�t�]i����FD�˥hS��P�W�h/ӊ����\�5B.���Ճk�f�o��K{��m���"�(HjI 